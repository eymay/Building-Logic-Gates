* NGSPICE file created from NOR2_eymenunay_pex.ext - technology: sky130B

.subckt NOR2_eymenunay_pex IN1 IN2 DVDD DGND OUT
X0 OUT.t1 IN2.t0 a_676_n108.t0 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 OUT.t0 IN2.t1 DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_676_n108.t1 IN1.t0 DVDD.t2 DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 OUT.t2 IN1.t1 DGND.t3 DGND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 IN2.n0 IN2.t0 248.348
R1 IN2.n0 IN2.t1 233.883
R2 IN2.n1 IN2.n0 0.542
R3 IN2 IN2.n1 0.062
R4 IN2.n1 IN2 0.062
R5 a_676_n108.t0 a_676_n108.t1 57.696
R6 OUT OUT.t1 29.863
R7 OUT.n0 OUT.t2 20.425
R8 OUT.n0 OUT.t0 18.375
R9 OUT OUT.n0 0.432
R10 DVDD.n18 DVDD.n14 497.647
R11 DVDD.n19 DVDD.n13 497.647
R12 DVDD.n11 DVDD.n7 140.046
R13 DVDD.n21 DVDD.n20 99.387
R14 DVDD.n16 DVDD.n15 53.082
R15 DVDD.n20 DVDD.n12 53.082
R16 DVDD.n12 DVDD.n11 53.082
R17 DVDD.n17 DVDD.n16 53.082
R18 DVDD.n26 DVDD.t2 28.859
R19 DVDD DVDD.n26 0.285
R20 DVDD.n23 DVDD.n22 0.167
R21 DVDD.n22 DVDD.n21 0.167
R22 DVDD.n4 DVDD.n1 0.109
R23 DVDD.n1 DVDD.n0 0.109
R24 DVDD.t0 DVDD.n8 0.034
R25 DVDD.n20 DVDD.n19 0.034
R26 DVDD.n19 DVDD.t1 0.034
R27 DVDD.n11 DVDD.n10 0.034
R28 DVDD.t1 DVDD.n18 0.034
R29 DVDD.n18 DVDD.n17 0.034
R30 DVDD.n4 DVDD.n3 0.031
R31 DVDD.n3 DVDD.n2 0.031
R32 DVDD.n10 DVDD.n9 0.029
R33 DVDD.n7 DVDD.n6 0.016
R34 DVDD.n24 DVDD.n23 0.006
R35 DVDD.n9 DVDD.t0 0.006
R36 DVDD.n25 DVDD.n24 0.006
R37 DVDD.n26 DVDD.n25 0.003
R38 DVDD.n5 DVDD.n4 0.001
R39 DVDD.n23 DVDD.n5 0.001
R40 DGND.n4 DGND.n1 816.97
R41 DGND.n23 DGND.n20 538.852
R42 DGND.n10 DGND.n9 138.164
R43 DGND.n8 DGND.n5 103.905
R44 DGND.n32 DGND.n29 93.74
R45 DGND.n5 DGND.n0 53.082
R46 DGND.n22 DGND.n21 35.011
R47 DGND.n33 DGND.n32 34.635
R48 DGND.n15 DGND.n8 34.258
R49 DGND.n22 DGND.t1 17.98
R50 DGND.n3 DGND.n2 17.898
R51 DGND.n28 DGND.n27 17.898
R52 DGND.n13 DGND.n12 17.789
R53 DGND.t0 DGND.t2 17.789
R54 DGND.n34 DGND.t3 17.689
R55 DGND.n16 DGND.t0 11.859
R56 DGND.n33 DGND.n15 9.788
R57 DGND.n32 DGND.n31 1.081
R58 DGND.n31 DGND.n30 1.081
R59 DGND.n26 DGND.n25 0.443
R60 DGND.n27 DGND.n26 0.443
R61 DGND.n8 DGND.n7 0.351
R62 DGND.n7 DGND.n6 0.351
R63 DGND DGND.n34 0.305
R64 DGND.n24 DGND.n19 0.218
R65 DGND.n19 DGND.n18 0.218
R66 DGND.n5 DGND.n4 0.109
R67 DGND.n4 DGND.n3 0.109
R68 DGND.n29 DGND.n28 0.109
R69 DGND.n15 DGND.n14 0.104
R70 DGND.n14 DGND.n13 0.104
R71 DGND.n11 DGND.n10 0.052
R72 DGND.n12 DGND.n11 0.052
R73 DGND.n24 DGND.n23 0.014
R74 DGND.n23 DGND.n22 0.014
R75 DGND.n33 DGND.n17 0.004
R76 DGND.n17 DGND.n16 0.004
R77 DGND.n34 DGND.n33 0.002
R78 DGND.n27 DGND.n24 0.001
R79 IN1.n0 IN1.t0 248.356
R80 IN1.n0 IN1.t1 233.881
R81 IN1 IN1.n0 0.648
C0 DVDD OUT 0.17fF
C1 IN2 OUT 0.25fF
C2 DVDD IN2 0.14fF
C3 IN1 OUT 0.02fF
C4 DVDD IN1 0.27fF
C5 IN1 IN2 0.07fF
.ends

