** sch_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/NOR2_eymenunay_TB.sch
**.subckt NOR2_eymenunay_TB
VDD VDD GND 1.8
V2 IN1 GND pulse 0 1.8 50n 1n 1n 100n 200n
V1 IN2 GND pulse 0 1.8 0n 1n 1n 100n 200n
X1 IN1 IN2 VDD GND OUT NOR2_eymenunay
C1 OUT GND 100f m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm




.control

tran 0.1n 400n
save all
plot  OUT

write NAND2_eymenunay.raw

.endc


**** end user architecture code
**.ends

* expanding   symbol:  NOR2_eymenunay.sym # of pins=5
** sym_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/NOR2_eymenunay.sym
** sch_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/NOR2_eymenunay.sch
.subckt NOR2_eymenunay  IN1 IN2 DVDD DGND OUT
*.ipin IN1
*.ipin IN2
*.opin OUT
*.iopin DVDD
*.iopin DGND
XM1 OUT IN1 DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN2 DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 IN1 DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT IN2 net1 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
