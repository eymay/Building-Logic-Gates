magic
tech sky130B
magscale 1 2
timestamp 1679245019
<< nwell >>
rect 450 -328 1192 240
<< pwell >>
rect 770 -354 1192 -351
rect 450 -909 1192 -354
rect 450 -912 872 -909
<< nmos >>
rect 646 -764 676 -564
rect 966 -761 996 -561
<< pmos >>
rect 646 -108 676 92
rect 966 -108 996 92
<< ndiff >>
rect 588 -576 646 -564
rect 588 -752 600 -576
rect 634 -752 646 -576
rect 588 -764 646 -752
rect 676 -576 734 -564
rect 676 -752 688 -576
rect 722 -752 734 -576
rect 676 -764 734 -752
rect 908 -573 966 -561
rect 908 -749 920 -573
rect 954 -749 966 -573
rect 908 -761 966 -749
rect 996 -573 1054 -561
rect 996 -749 1008 -573
rect 1042 -749 1054 -573
rect 996 -761 1054 -749
<< pdiff >>
rect 588 80 646 92
rect 588 -96 600 80
rect 634 -96 646 80
rect 588 -108 646 -96
rect 676 80 734 92
rect 676 -96 688 80
rect 722 -96 734 80
rect 676 -108 734 -96
rect 908 80 966 92
rect 908 -96 920 80
rect 954 -96 966 80
rect 908 -108 966 -96
rect 996 80 1054 92
rect 996 -96 1008 80
rect 1042 -96 1054 80
rect 996 -108 1054 -96
<< ndiffc >>
rect 600 -752 634 -576
rect 688 -752 722 -576
rect 920 -749 954 -573
rect 1008 -749 1042 -573
<< pdiffc >>
rect 600 -96 634 80
rect 688 -96 722 80
rect 920 -96 954 80
rect 1008 -96 1042 80
<< psubdiff >>
rect 806 -390 902 -387
rect 486 -424 582 -390
rect 740 -421 902 -390
rect 1060 -421 1156 -387
rect 740 -424 840 -421
rect 486 -486 520 -424
rect 486 -842 520 -780
rect 802 -839 840 -424
rect 1122 -483 1156 -421
rect 1122 -839 1156 -777
rect 802 -842 902 -839
rect 486 -876 582 -842
rect 740 -873 902 -842
rect 1060 -873 1156 -839
rect 740 -876 836 -873
<< nsubdiff >>
rect 486 170 582 204
rect 740 170 902 204
rect 1060 170 1156 204
rect 486 107 520 170
rect 486 -258 520 -195
rect 802 -258 840 170
rect 1122 107 1156 170
rect 1122 -258 1156 -195
rect 486 -292 582 -258
rect 740 -292 902 -258
rect 1060 -292 1156 -258
<< psubdiffcont >>
rect 582 -424 740 -390
rect 902 -421 1060 -387
rect 486 -780 520 -486
rect 1122 -777 1156 -483
rect 582 -876 740 -842
rect 902 -873 1060 -839
<< nsubdiffcont >>
rect 582 170 740 204
rect 902 170 1060 204
rect 486 -195 520 107
rect 1122 -195 1156 107
rect 582 -292 740 -258
rect 902 -292 1060 -258
<< poly >>
rect 646 92 676 118
rect 646 -139 676 -108
rect 628 -155 694 -139
rect 628 -189 644 -155
rect 678 -189 694 -155
rect 628 -205 694 -189
rect 966 92 996 118
rect 966 -139 996 -108
rect 948 -155 1014 -139
rect 948 -189 964 -155
rect 998 -189 1014 -155
rect 948 -205 1014 -189
rect 628 -492 694 -476
rect 628 -526 644 -492
rect 678 -526 694 -492
rect 628 -542 694 -526
rect 646 -564 676 -542
rect 646 -790 676 -764
rect 948 -489 1014 -473
rect 948 -523 964 -489
rect 998 -523 1014 -489
rect 948 -539 1014 -523
rect 966 -561 996 -539
rect 966 -787 996 -761
<< polycont >>
rect 644 -189 678 -155
rect 964 -189 998 -155
rect 644 -526 678 -492
rect 964 -523 998 -489
<< locali >>
rect 486 170 582 204
rect 740 170 902 204
rect 1060 170 1156 204
rect 486 107 520 170
rect 600 80 634 96
rect 600 -112 634 -96
rect 688 80 722 96
rect 688 -112 722 -96
rect 628 -189 644 -155
rect 678 -189 694 -155
rect 486 -258 520 -195
rect 802 -258 840 170
rect 1122 107 1156 170
rect 920 80 954 96
rect 920 -112 954 -96
rect 1008 80 1042 96
rect 1008 -112 1042 -96
rect 948 -189 964 -155
rect 998 -189 1014 -155
rect 1122 -258 1156 -195
rect 486 -292 582 -258
rect 740 -292 902 -258
rect 1060 -292 1156 -258
rect 806 -390 902 -387
rect 486 -424 582 -390
rect 740 -421 902 -390
rect 1060 -421 1156 -387
rect 740 -424 840 -421
rect 486 -486 520 -424
rect 628 -526 644 -492
rect 678 -526 694 -492
rect 600 -576 634 -560
rect 600 -768 634 -752
rect 688 -576 722 -560
rect 688 -768 722 -752
rect 486 -842 520 -780
rect 802 -839 840 -424
rect 1122 -483 1156 -421
rect 948 -523 964 -489
rect 998 -523 1014 -489
rect 920 -573 954 -557
rect 920 -765 954 -749
rect 1008 -573 1042 -557
rect 1008 -765 1042 -749
rect 1122 -839 1156 -777
rect 802 -842 902 -839
rect 486 -876 582 -842
rect 740 -873 902 -842
rect 1060 -873 1156 -839
rect 740 -876 836 -873
<< viali >>
rect 486 -83 520 22
rect 600 -96 634 80
rect 688 -96 722 80
rect 644 -189 678 -155
rect 920 -96 954 80
rect 1008 -96 1042 80
rect 964 -189 998 -155
rect 644 -526 678 -492
rect 486 -721 520 -597
rect 600 -752 634 -576
rect 688 -752 722 -576
rect 964 -523 998 -489
rect 920 -749 954 -573
rect 1008 -749 1042 -573
rect 902 -873 965 -839
<< metal1 >>
rect 594 80 640 92
rect 235 -16 435 65
rect 480 22 526 34
rect 480 -16 486 22
rect 235 -69 486 -16
rect 235 -135 435 -69
rect 480 -83 486 -69
rect 520 -16 526 22
rect 594 -16 600 80
rect 520 -69 600 -16
rect 520 -83 526 -69
rect 480 -95 526 -83
rect 594 -96 600 -69
rect 634 -96 640 80
rect 594 -108 640 -96
rect 682 80 728 92
rect 682 -96 688 80
rect 722 2 728 80
rect 914 80 960 92
rect 914 2 920 80
rect 722 -50 920 2
rect 722 -96 728 -50
rect 682 -108 728 -96
rect 914 -96 920 -50
rect 954 -96 960 80
rect 914 -108 960 -96
rect 1002 80 1048 92
rect 1002 -96 1008 80
rect 1042 8 1048 80
rect 1042 -48 1402 8
rect 1042 -96 1048 -48
rect 1002 -108 1048 -96
rect 632 -155 690 -149
rect 632 -189 644 -155
rect 678 -189 690 -155
rect 235 -320 435 -242
rect 632 -320 690 -189
rect 235 -367 690 -320
rect 235 -442 435 -367
rect 632 -492 690 -367
rect 632 -526 644 -492
rect 678 -526 690 -492
rect 632 -532 690 -526
rect 952 -155 1010 -149
rect 952 -189 964 -155
rect 998 -189 1010 -155
rect 952 -316 1010 -189
rect 1345 -224 1401 -48
rect 1214 -316 1306 -294
rect 952 -363 1306 -316
rect 952 -489 1010 -363
rect 1214 -386 1306 -363
rect 1336 -424 1536 -224
rect 952 -523 964 -489
rect 998 -523 1010 -489
rect 952 -529 1010 -523
rect 231 -640 431 -554
rect 594 -576 640 -564
rect 480 -597 526 -585
rect 480 -640 486 -597
rect 231 -690 486 -640
rect 231 -754 431 -690
rect 480 -721 486 -690
rect 520 -640 526 -597
rect 594 -640 600 -576
rect 520 -690 600 -640
rect 520 -721 526 -690
rect 480 -733 526 -721
rect 594 -752 600 -690
rect 634 -752 640 -576
rect 594 -764 640 -752
rect 682 -576 728 -564
rect 682 -752 688 -576
rect 722 -752 728 -576
rect 682 -764 728 -752
rect 914 -573 960 -561
rect 914 -749 920 -573
rect 954 -749 960 -573
rect 914 -761 960 -749
rect 1002 -573 1048 -561
rect 1002 -749 1008 -573
rect 1042 -579 1048 -573
rect 1371 -579 1423 -424
rect 1042 -628 1423 -579
rect 1042 -749 1048 -628
rect 1002 -761 1048 -749
rect 685 -919 722 -764
rect 921 -833 955 -761
rect 890 -839 977 -833
rect 890 -873 902 -839
rect 965 -873 977 -839
rect 890 -879 977 -873
rect 1371 -919 1423 -628
rect 685 -978 1427 -919
<< labels >>
flabel metal1 1214 -386 1306 -294 1 FreeMono 160 0 0 0 IN2
port 5 n
flabel metal1 1336 -424 1536 -224 0 FreeSans 256 0 0 0 OUT
port 4 nsew
flabel metal1 235 -442 435 -242 0 FreeSans 256 0 0 0 IN1
port 0 nsew
flabel metal1 231 -754 431 -554 0 FreeSans 256 0 0 0 DGND
port 3 nsew
flabel metal1 235 -135 435 65 0 FreeSans 256 0 0 0 DVDD
port 2 nsew
<< end >>
