magic
tech sky130B
magscale 1 2
timestamp 1679300852
<< locali >>
rect 1968 682 2002 870
rect 1963 215 1997 403
<< viali >>
rect 1091 1192 1128 1279
rect 1967 1020 2001 1088
rect 1089 714 1125 791
rect 1089 233 1125 310
rect 1783 -101 1866 -63
<< metal1 >>
rect 819 1271 1019 1385
rect 1570 1324 1770 1449
rect 1085 1279 1134 1291
rect 1085 1271 1091 1279
rect 819 1204 1091 1271
rect 819 1185 1019 1204
rect 1085 1192 1091 1204
rect 1128 1246 1134 1279
rect 1562 1254 1572 1324
rect 1625 1254 1770 1324
rect 1809 1258 2009 1458
rect 1570 1249 1770 1254
rect 1128 1197 1242 1246
rect 1128 1192 1134 1197
rect 1085 1180 1134 1192
rect 1285 1156 1295 1226
rect 1348 1156 1358 1226
rect 815 1023 1015 1095
rect 1710 1038 1761 1249
rect 1967 1100 2002 1258
rect 1961 1088 2007 1100
rect 1239 1023 1655 1025
rect 815 986 1655 1023
rect 1961 1020 1967 1088
rect 2001 1020 2007 1088
rect 1961 1008 2007 1020
rect 815 895 1015 986
rect 1239 982 1655 986
rect 1083 791 1131 803
rect 1083 714 1089 791
rect 1125 762 1131 791
rect 1125 715 1235 762
rect 1125 714 1131 715
rect 1083 702 1131 714
rect 1283 694 1293 764
rect 1346 694 1356 764
rect 809 563 1009 601
rect 1778 573 1836 984
rect 1236 563 1658 565
rect 809 526 1658 563
rect 809 401 1009 526
rect 1236 522 1658 526
rect 1083 310 1131 322
rect 1083 233 1089 310
rect 1125 280 1131 310
rect 1125 233 1232 280
rect 1083 221 1131 233
rect 1282 221 1292 291
rect 1345 221 1355 291
rect 825 101 1025 194
rect 1770 107 1828 518
rect 1235 101 1653 106
rect 825 64 1653 101
rect 825 -6 1025 64
rect 1783 -57 1846 44
rect 1771 -63 1878 -57
rect 1771 -101 1783 -63
rect 1866 -101 1878 -63
rect 1771 -107 1878 -101
<< via1 >>
rect 1572 1254 1625 1324
rect 1295 1156 1348 1226
rect 1293 694 1346 764
rect 1292 221 1345 291
<< metal2 >>
rect 1295 1318 1353 1328
rect 1572 1324 1625 1334
rect 1295 1254 1572 1318
rect 1295 1253 1625 1254
rect 1295 1226 1353 1253
rect 1572 1244 1625 1253
rect 1348 1156 1353 1226
rect 1295 774 1353 1156
rect 1293 764 1353 774
rect 1346 694 1353 764
rect 1293 684 1353 694
rect 1295 301 1353 684
rect 1292 291 1353 301
rect 1345 222 1353 291
rect 1292 211 1345 221
use sky130_fd_pr__nfet_01v8_64Z3AY  XM1
timestamp 1679299220
transform 0 -1 1754 1 0 76
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1679299220
transform 0 -1 1758 1 0 1009
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_QDT3BL  XM3
timestamp 1679299220
transform 1 0 1263 0 1 210
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_BDT3BC  XM4
timestamp 1679299220
transform 1 0 1265 0 1 672
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_7HS3BC  XM5
timestamp 1679299220
transform 1 0 1267 0 1 1132
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM6
timestamp 1679299220
transform 0 -1 1759 1 0 544
box -211 -279 211 279
<< labels >>
flabel metal1 809 401 1009 601 0 FreeSans 256 0 0 0 IN2
port 1 nsew
flabel metal1 819 1185 1019 1385 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal1 1809 1258 2009 1458 0 FreeSans 256 0 0 0 DGND
port 4 nsew
flabel metal1 1570 1249 1770 1449 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 825 -6 1025 194 0 FreeSans 256 0 0 0 IN3
port 5 nsew
flabel metal1 815 895 1015 1095 0 FreeSans 256 0 0 0 IN1
port 0 nsew
<< end >>
