magic
tech sky130B
magscale 1 2
timestamp 1679299220
<< error_s >>
rect 298 1097 333 1131
rect 299 1078 333 1097
rect 685 1078 738 1079
rect 129 1029 187 1035
rect 129 995 141 1029
rect 129 989 187 995
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 1078
rect 352 1044 387 1078
rect 667 1044 738 1078
rect 352 583 386 1044
rect 668 1043 738 1044
rect 685 1009 756 1043
rect 1036 1009 1071 1043
rect 498 976 556 982
rect 498 942 510 976
rect 498 936 556 942
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 685 530 755 1009
rect 1037 990 1071 1009
rect 867 941 925 947
rect 867 907 879 941
rect 867 901 925 907
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1056 477 1071 990
rect 1090 956 1125 990
rect 1405 956 1440 990
rect 1090 477 1124 956
rect 1406 937 1440 956
rect 1236 888 1294 894
rect 1236 854 1248 888
rect 1236 848 1294 854
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 937
rect 1459 903 1494 937
rect 1774 903 1809 920
rect 1459 424 1493 903
rect 1775 902 1809 903
rect 1775 866 1845 902
rect 1605 835 1663 841
rect 1605 801 1617 835
rect 1792 832 1863 866
rect 1605 795 1663 801
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 832
rect 1974 764 2032 770
rect 1974 730 1986 764
rect 1974 724 2032 730
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1679299220
transform 1 0 158 0 1 857
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1679299220
transform 1 0 527 0 1 804
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1679299220
transform 1 0 896 0 1 760
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1679299220
transform 1 0 1265 0 1 707
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM5
timestamp 1679299220
transform 1 0 1634 0 1 654
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1679299220
transform 1 0 2003 0 1 592
box -211 -310 211 310
<< end >>
