* NGSPICE file created from NAND3_eymenunay_pex.ext - technology: sky130B

.subckt NAND3_eymenunay_pex IN1 IN2 OUT IN3 DVDD DGND
X0 OUT IN3.t0 DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=150000u
X1 a_1685_91.t0 IN3.t1 DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 OUT.t1 IN1.t0 DVDD.t3 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 OUT.t3 IN1.t1 a_1689_936.t0 DGND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 OUT IN2.t0 DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1689_936.t1 IN2.t1 a_1685_91.t1 DGND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 IN3.n0 IN3.t0 247.986
R1 IN3.n0 IN3.t1 234.588
R2 IN3 IN3.n0 0.907
R3 DVDD.n1 DVDD.n0 762.352
R4 DVDD.n46 DVDD.n45 754.901
R5 DVDD.n20 DVDD.n7 321.175
R6 DVDD.n30 DVDD.n29 278.43
R7 DVDD.t2 DVDD.t4 241.981
R8 DVDD.n50 DVDD.n47 140.046
R9 DVDD.n22 DVDD.n6 118.211
R10 DVDD.n11 DVDD.n10 115.952
R11 DVDD.n35 DVDD.n3 111.644
R12 DVDD.n31 DVDD.n30 94.722
R13 DVDD.n43 DVDD.n42 86.467
R14 DVDD.n51 DVDD.n50 83.952
R15 DVDD.n6 DVDD.n5 80.564
R16 DVDD.n3 DVDD.n2 79.811
R17 DVDD.n36 DVDD.n35 62.494
R18 DVDD.n23 DVDD.n22 59.858
R19 DVDD.n22 DVDD.n21 34.257
R20 DVDD.n35 DVDD.n34 29.699
R21 DVDD.n52 DVDD.t3 28.901
R22 DVDD.n33 DVDD.t5 28.857
R23 DVDD.n17 DVDD.t1 28.832
R24 DVDD.n34 DVDD.n33 19.889
R25 DVDD.n52 DVDD.n51 15.973
R26 DVDD.n18 DVDD.n17 8.855
R27 DVDD.n19 DVDD.n18 8.567
R28 DVDD.n21 DVDD.n20 0.502
R29 DVDD.n20 DVDD.n19 0.482
R30 DVDD DVDD.n52 0.274
R31 DVDD.n15 DVDD.n12 0.061
R32 DVDD.n12 DVDD.n11 0.061
R33 DVDD.n27 DVDD.n24 0.053
R34 DVDD.n24 DVDD.n23 0.053
R35 DVDD.n40 DVDD.n37 0.048
R36 DVDD.n37 DVDD.n36 0.048
R37 DVDD.n50 DVDD.n49 0.034
R38 DVDD.n10 DVDD.n9 0.034
R39 DVDD.n15 DVDD.n14 0.031
R40 DVDD.n27 DVDD.n26 0.031
R41 DVDD.n40 DVDD.n39 0.031
R42 DVDD.n26 DVDD.n25 0.031
R43 DVDD.n14 DVDD.n13 0.031
R44 DVDD.n39 DVDD.n38 0.031
R45 DVDD.n49 DVDD.n48 0.028
R46 DVDD.n9 DVDD.n8 0.028
R47 DVDD.n19 DVDD.n16 0.02
R48 DVDD.n47 DVDD.n46 0.016
R49 DVDD.n5 DVDD.n4 0.016
R50 DVDD.n2 DVDD.n1 0.016
R51 DVDD.n33 DVDD.n32 0.01
R52 DVDD.n52 DVDD.n44 0.008
R53 DVDD.n48 DVDD.t2 0.007
R54 DVDD.n8 DVDD.t0 0.007
R55 DVDD.n32 DVDD.n31 0.006
R56 DVDD.n31 DVDD.n28 0.005
R57 DVDD.n43 DVDD.n41 0.005
R58 DVDD.n44 DVDD.n43 0.004
R59 DVDD.n41 DVDD.n40 0.001
R60 DVDD.n28 DVDD.n27 0.001
R61 DVDD.n16 DVDD.n15 0.001
R62 OUT.n0 OUT.t1 29.272
R63 OUT.n0 OUT.t3 18.045
R64 OUT OUT.n0 0.017
R65 DGND.n3 DGND.t3 323.222
R66 DGND.n36 DGND.t2 323.222
R67 DGND.n26 DGND.t0 323.222
R68 DGND.n7 DGND.n6 138.164
R69 DGND.n28 DGND.n14 138.164
R70 DGND.n39 DGND.n33 138.164
R71 DGND.n47 DGND.n7 121.223
R72 DGND.n29 DGND.n28 85.082
R73 DGND.n40 DGND.n39 85.082
R74 DGND.n31 DGND.n30 54.964
R75 DGND.n40 DGND.n31 53.082
R76 DGND.n29 DGND.n12 53.082
R77 DGND.n41 DGND.n40 49.511
R78 DGND.n42 DGND.n41 46.477
R79 DGND.n30 DGND.n29 44.423
R80 DGND.n17 DGND.n16 26.59
R81 DGND.n24 DGND.n20 24.727
R82 DGND.n24 DGND.n23 22.211
R83 DGND.n20 DGND.n17 20.547
R84 DGND.n20 DGND.t1 17.63
R85 DGND.n16 DGND.n15 15.171
R86 DGND DGND.n47 0.804
R87 DGND.n43 DGND.n42 0.482
R88 DGND.n44 DGND.n43 0.481
R89 DGND.n9 DGND.n8 0.218
R90 DGND.n44 DGND.n9 0.218
R91 DGND.n23 DGND.n22 0.19
R92 DGND.n6 DGND.n5 0.109
R93 DGND.n31 DGND.n10 0.109
R94 DGND.n12 DGND.n11 0.109
R95 DGND.n14 DGND.n13 0.109
R96 DGND.n33 DGND.n32 0.109
R97 DGND.n25 DGND.n24 0.104
R98 DGND.n26 DGND.n25 0.104
R99 DGND.n22 DGND.n21 0.097
R100 DGND.n7 DGND.n4 0.052
R101 DGND.n4 DGND.n3 0.052
R102 DGND.n1 DGND.n0 0.052
R103 DGND.n28 DGND.n27 0.052
R104 DGND.n27 DGND.n26 0.052
R105 DGND.n35 DGND.n34 0.052
R106 DGND.n36 DGND.n35 0.052
R107 DGND.n39 DGND.n38 0.052
R108 DGND.n3 DGND.n2 0.028
R109 DGND.n37 DGND.n36 0.028
R110 DGND.n2 DGND.n1 0.025
R111 DGND.n38 DGND.n37 0.025
R112 DGND.n47 DGND.n46 0.012
R113 DGND.n46 DGND.n45 0.012
R114 DGND.n20 DGND.n19 0.008
R115 DGND.n19 DGND.n18 0.008
R116 DGND.n45 DGND.n44 0.001
R117 a_1685_91.t0 a_1685_91.t1 35.627
R118 IN1.n0 IN1.t0 247.986
R119 IN1.n0 IN1.t1 234.568
R120 IN1 IN1.n0 0.956
R121 a_1689_936.t0 a_1689_936.t1 35.621
R122 IN2.n0 IN2.t0 247.986
R123 IN2.n0 IN2.t1 234.577
R124 IN2 IN2.n0 0.969
C0 IN3 IN1 0.01fF
C1 IN3 IN2 0.09fF
C2 OUT IN1 0.14fF
C3 IN2 OUT 0.10fF
C4 IN1 DVDD 0.42fF
C5 IN2 DVDD 0.35fF
C6 IN3 OUT 0.09fF
C7 IN3 DVDD 0.30fF
C8 OUT DVDD 1.32fF
C9 IN2 IN1 0.08fF
.ends

