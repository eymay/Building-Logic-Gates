magic
tech sky130B
magscale 1 2
timestamp 1679301765
<< nwell >>
rect 1056 956 1478 1416
rect 1054 848 1478 956
rect 1054 494 1476 848
rect 1052 388 1476 494
rect 1052 -74 1474 388
<< pwell >>
rect 1479 798 2037 1220
rect 1480 333 2038 755
rect 1475 -135 2033 287
<< nmos >>
rect 1689 994 1889 1024
rect 1690 529 1890 559
rect 1685 61 1885 91
<< pmos >>
rect 1252 1068 1282 1268
rect 1250 608 1280 808
rect 1248 146 1278 346
<< ndiff >>
rect 1689 1070 1889 1082
rect 1689 1036 1701 1070
rect 1877 1036 1889 1070
rect 1689 1024 1889 1036
rect 1689 982 1889 994
rect 1689 948 1701 982
rect 1877 948 1889 982
rect 1689 936 1889 948
rect 1690 605 1890 617
rect 1690 571 1702 605
rect 1878 571 1890 605
rect 1690 559 1890 571
rect 1690 517 1890 529
rect 1690 483 1702 517
rect 1878 483 1890 517
rect 1690 471 1890 483
rect 1685 137 1885 149
rect 1685 103 1697 137
rect 1873 103 1885 137
rect 1685 91 1885 103
rect 1685 49 1885 61
rect 1685 15 1697 49
rect 1873 15 1885 49
rect 1685 3 1885 15
<< pdiff >>
rect 1194 1256 1252 1268
rect 1194 1080 1206 1256
rect 1240 1080 1252 1256
rect 1194 1068 1252 1080
rect 1282 1256 1340 1268
rect 1282 1080 1294 1256
rect 1328 1080 1340 1256
rect 1282 1068 1340 1080
rect 1192 796 1250 808
rect 1192 620 1204 796
rect 1238 620 1250 796
rect 1192 608 1250 620
rect 1280 796 1338 808
rect 1280 620 1292 796
rect 1326 620 1338 796
rect 1280 608 1338 620
rect 1190 334 1248 346
rect 1190 158 1202 334
rect 1236 158 1248 334
rect 1190 146 1248 158
rect 1278 334 1336 346
rect 1278 158 1290 334
rect 1324 158 1336 334
rect 1278 146 1336 158
<< ndiffc >>
rect 1701 1036 1877 1070
rect 1701 948 1877 982
rect 1702 571 1878 605
rect 1702 483 1878 517
rect 1697 103 1873 137
rect 1697 15 1873 49
<< pdiffc >>
rect 1206 1080 1240 1256
rect 1294 1080 1328 1256
rect 1204 620 1238 796
rect 1292 620 1326 796
rect 1202 158 1236 334
rect 1290 158 1324 334
<< psubdiff >>
rect 1515 1150 1611 1184
rect 1905 1150 2001 1184
rect 1515 1088 1549 1150
rect 1967 1088 2001 1150
rect 1515 868 1549 930
rect 1967 868 2001 930
rect 1515 834 1611 868
rect 1905 834 2001 868
rect 1516 685 1612 719
rect 1906 685 2002 719
rect 1516 623 1550 685
rect 1968 623 2002 685
rect 1516 403 1550 465
rect 1968 403 2002 465
rect 1516 369 1612 403
rect 1906 369 2002 403
rect 1511 217 1607 251
rect 1901 217 1997 251
rect 1511 155 1545 217
rect 1963 155 1997 217
rect 1511 -65 1545 -3
rect 1963 -65 1997 -3
rect 1511 -99 1607 -65
rect 1901 -99 1997 -65
<< nsubdiff >>
rect 1092 1346 1188 1380
rect 1346 1346 1442 1380
rect 1092 1283 1126 1346
rect 1408 1283 1442 1346
rect 1092 920 1126 981
rect 1408 920 1442 981
rect 1090 884 1442 920
rect 1090 823 1124 884
rect 1406 823 1440 884
rect 1090 458 1124 521
rect 1406 458 1440 521
rect 1088 424 1440 458
rect 1088 361 1122 424
rect 1404 361 1438 424
rect 1088 -4 1122 59
rect 1404 -4 1438 59
rect 1088 -38 1184 -4
rect 1342 -38 1438 -4
<< psubdiffcont >>
rect 1611 1150 1905 1184
rect 1515 930 1549 1088
rect 1967 930 2001 1088
rect 1611 834 1905 868
rect 1612 685 1906 719
rect 1516 465 1550 623
rect 1968 465 2002 623
rect 1612 369 1906 403
rect 1607 217 1901 251
rect 1511 -3 1545 155
rect 1963 -3 1997 155
rect 1607 -99 1901 -65
<< nsubdiffcont >>
rect 1188 1346 1346 1380
rect 1092 981 1126 1283
rect 1408 981 1442 1283
rect 1090 521 1124 823
rect 1406 521 1440 823
rect 1088 59 1122 361
rect 1404 59 1438 361
rect 1184 -38 1342 -4
<< poly >>
rect 1252 1268 1282 1294
rect 1252 1037 1282 1068
rect 1234 1021 1300 1037
rect 1234 987 1250 1021
rect 1284 987 1300 1021
rect 1234 971 1300 987
rect 1601 1026 1667 1042
rect 1601 992 1617 1026
rect 1651 1024 1667 1026
rect 1651 994 1689 1024
rect 1889 994 1915 1024
rect 1651 992 1667 994
rect 1601 976 1667 992
rect 1250 808 1280 834
rect 1250 577 1280 608
rect 1232 561 1298 577
rect 1232 527 1248 561
rect 1282 527 1298 561
rect 1232 511 1298 527
rect 1602 561 1668 577
rect 1602 527 1618 561
rect 1652 559 1668 561
rect 1652 529 1690 559
rect 1890 529 1916 559
rect 1652 527 1668 529
rect 1602 511 1668 527
rect 1248 346 1278 372
rect 1248 115 1278 146
rect 1230 99 1296 115
rect 1230 65 1246 99
rect 1280 65 1296 99
rect 1230 49 1296 65
rect 1597 93 1663 109
rect 1597 59 1613 93
rect 1647 91 1663 93
rect 1647 61 1685 91
rect 1885 61 1911 91
rect 1647 59 1663 61
rect 1597 43 1663 59
<< polycont >>
rect 1250 987 1284 1021
rect 1617 992 1651 1026
rect 1248 527 1282 561
rect 1618 527 1652 561
rect 1246 65 1280 99
rect 1613 59 1647 93
<< locali >>
rect 1092 1346 1188 1380
rect 1346 1346 1442 1380
rect 1092 1283 1126 1346
rect 1408 1283 1442 1346
rect 1206 1256 1240 1272
rect 1206 1064 1240 1080
rect 1294 1256 1328 1272
rect 1294 1064 1328 1080
rect 1234 987 1250 1021
rect 1284 987 1300 1021
rect 1092 920 1126 981
rect 1408 920 1442 981
rect 1090 884 1442 920
rect 1515 1150 1611 1184
rect 1905 1150 2001 1184
rect 1515 1088 1549 1150
rect 1967 1088 2001 1150
rect 1617 1026 1651 1042
rect 1685 1036 1701 1070
rect 1877 1036 1893 1070
rect 1617 976 1651 992
rect 1685 948 1701 982
rect 1877 948 1893 982
rect 1090 823 1124 884
rect 1406 823 1440 884
rect 1515 868 1549 930
rect 1967 870 2001 930
rect 1967 868 2002 870
rect 1515 834 1611 868
rect 1905 834 2002 868
rect 1204 796 1238 812
rect 1204 604 1238 620
rect 1292 796 1326 812
rect 1292 604 1326 620
rect 1232 527 1248 561
rect 1282 527 1298 561
rect 1090 458 1124 521
rect 1968 719 2002 834
rect 1406 458 1440 521
rect 1088 424 1440 458
rect 1516 685 1612 719
rect 1906 685 2002 719
rect 1516 623 1550 685
rect 1968 623 2002 685
rect 1618 561 1652 577
rect 1686 571 1702 605
rect 1878 571 1894 605
rect 1618 511 1652 527
rect 1686 483 1702 517
rect 1878 483 1894 517
rect 1088 361 1122 424
rect 1404 361 1438 424
rect 1516 403 1550 465
rect 1968 403 2002 465
rect 1516 369 1612 403
rect 1906 369 2002 403
rect 1202 334 1236 350
rect 1202 142 1236 158
rect 1290 334 1324 350
rect 1290 142 1324 158
rect 1230 65 1246 99
rect 1280 65 1296 99
rect 1088 -4 1122 59
rect 1963 251 1997 369
rect 1404 -4 1438 59
rect 1088 -38 1184 -4
rect 1342 -38 1438 -4
rect 1511 217 1607 251
rect 1901 217 1997 251
rect 1511 155 1545 217
rect 1963 155 1997 217
rect 1613 93 1647 109
rect 1681 103 1697 137
rect 1873 103 1889 137
rect 1613 43 1647 59
rect 1681 15 1697 49
rect 1873 15 1889 49
rect 1511 -65 1545 -3
rect 1963 -65 1997 -3
rect 1511 -99 1607 -65
rect 1901 -99 1997 -65
<< viali >>
rect 1091 1192 1092 1279
rect 1092 1192 1126 1279
rect 1126 1192 1128 1279
rect 1206 1080 1240 1256
rect 1294 1080 1328 1256
rect 1250 987 1284 1021
rect 1701 1036 1877 1070
rect 1617 992 1651 1026
rect 1967 1020 2001 1088
rect 1701 948 1877 982
rect 1089 714 1090 791
rect 1090 714 1124 791
rect 1124 714 1125 791
rect 1204 620 1238 796
rect 1292 620 1326 796
rect 1248 527 1282 561
rect 1702 571 1878 605
rect 1618 527 1652 561
rect 1702 483 1878 517
rect 1089 233 1122 310
rect 1122 233 1125 310
rect 1202 158 1236 334
rect 1290 158 1324 334
rect 1246 65 1280 99
rect 1697 103 1873 137
rect 1613 59 1647 93
rect 1697 15 1873 49
rect 1783 -65 1866 -63
rect 1783 -99 1866 -65
rect 1783 -101 1866 -99
<< metal1 >>
rect 819 1271 1019 1385
rect 1570 1324 1770 1449
rect 1085 1279 1134 1291
rect 1085 1271 1091 1279
rect 819 1204 1091 1271
rect 819 1185 1019 1204
rect 1085 1192 1091 1204
rect 1128 1246 1134 1279
rect 1200 1256 1246 1268
rect 1200 1246 1206 1256
rect 1128 1197 1206 1246
rect 1128 1192 1134 1197
rect 1085 1180 1134 1192
rect 815 1023 1015 1095
rect 1200 1080 1206 1197
rect 1240 1080 1246 1256
rect 1288 1256 1334 1268
rect 1288 1226 1294 1256
rect 1328 1226 1334 1256
rect 1562 1254 1572 1324
rect 1625 1254 1770 1324
rect 1809 1258 2009 1458
rect 1570 1249 1770 1254
rect 1285 1156 1294 1226
rect 1348 1156 1358 1226
rect 1200 1068 1246 1080
rect 1288 1080 1294 1156
rect 1328 1080 1334 1156
rect 1288 1068 1334 1080
rect 1710 1076 1761 1249
rect 1967 1100 2002 1258
rect 1961 1088 2007 1100
rect 1689 1070 1889 1076
rect 1238 1025 1296 1027
rect 1611 1026 1657 1038
rect 1689 1036 1701 1070
rect 1877 1036 1889 1070
rect 1689 1030 1889 1036
rect 1611 1025 1617 1026
rect 1238 1023 1617 1025
rect 815 1021 1617 1023
rect 815 987 1250 1021
rect 1284 992 1617 1021
rect 1651 992 1657 1026
rect 1961 1020 1967 1088
rect 2001 1020 2007 1088
rect 1961 1008 2007 1020
rect 1284 987 1657 992
rect 815 986 1657 987
rect 815 895 1015 986
rect 1238 982 1657 986
rect 1238 981 1296 982
rect 1611 980 1657 982
rect 1689 982 1889 988
rect 1689 948 1701 982
rect 1877 948 1889 982
rect 1689 942 1889 948
rect 1083 791 1131 803
rect 1083 714 1089 791
rect 1125 762 1131 791
rect 1198 796 1244 808
rect 1198 762 1204 796
rect 1125 715 1204 762
rect 1125 714 1131 715
rect 1083 702 1131 714
rect 1198 620 1204 715
rect 1238 620 1244 796
rect 1286 796 1332 808
rect 1286 764 1292 796
rect 1326 764 1332 796
rect 1283 694 1292 764
rect 1346 694 1356 764
rect 1198 608 1244 620
rect 1286 620 1292 694
rect 1326 620 1332 694
rect 1286 608 1332 620
rect 1778 611 1836 942
rect 1690 605 1890 611
rect 809 563 1009 601
rect 1236 565 1294 567
rect 1612 565 1658 573
rect 1690 571 1702 605
rect 1878 571 1890 605
rect 1690 565 1890 571
rect 1236 563 1658 565
rect 809 561 1658 563
rect 809 527 1248 561
rect 1282 527 1618 561
rect 1652 527 1658 561
rect 809 526 1658 527
rect 809 401 1009 526
rect 1236 522 1658 526
rect 1236 521 1294 522
rect 1612 515 1658 522
rect 1690 517 1890 523
rect 1690 483 1702 517
rect 1878 483 1890 517
rect 1690 477 1890 483
rect 1196 334 1242 346
rect 1083 310 1131 322
rect 1083 233 1089 310
rect 1125 280 1131 310
rect 1196 280 1202 334
rect 1125 233 1202 280
rect 1083 221 1131 233
rect 825 101 1025 194
rect 1196 158 1202 233
rect 1236 158 1242 334
rect 1284 334 1330 346
rect 1284 291 1290 334
rect 1324 291 1330 334
rect 1282 221 1290 291
rect 1345 221 1355 291
rect 1196 146 1242 158
rect 1284 158 1290 221
rect 1324 158 1330 221
rect 1284 146 1330 158
rect 1770 143 1828 477
rect 1685 137 1885 143
rect 1235 105 1653 106
rect 1234 101 1653 105
rect 825 99 1653 101
rect 825 65 1246 99
rect 1280 93 1653 99
rect 1685 103 1697 137
rect 1873 103 1885 137
rect 1685 97 1885 103
rect 1280 65 1613 93
rect 825 64 1613 65
rect 825 -6 1025 64
rect 1234 59 1292 64
rect 1607 59 1613 64
rect 1647 59 1653 93
rect 1607 47 1653 59
rect 1685 49 1885 55
rect 1685 15 1697 49
rect 1873 15 1885 49
rect 1685 9 1885 15
rect 1783 -57 1846 9
rect 1771 -63 1878 -57
rect 1771 -101 1783 -63
rect 1866 -101 1878 -63
rect 1771 -107 1878 -101
<< via1 >>
rect 1572 1254 1625 1324
rect 1295 1156 1328 1226
rect 1328 1156 1348 1226
rect 1293 694 1326 764
rect 1326 694 1346 764
rect 1292 221 1324 291
rect 1324 221 1345 291
<< metal2 >>
rect 1295 1318 1353 1328
rect 1572 1324 1625 1334
rect 1295 1254 1572 1318
rect 1295 1253 1625 1254
rect 1295 1226 1353 1253
rect 1572 1244 1625 1253
rect 1348 1156 1353 1226
rect 1295 774 1353 1156
rect 1293 764 1353 774
rect 1346 694 1353 764
rect 1293 684 1353 694
rect 1295 301 1353 684
rect 1292 291 1353 301
rect 1345 222 1353 291
rect 1292 211 1345 221
<< labels >>
flabel metal1 809 401 1009 601 0 FreeSans 256 0 0 0 IN2
port 1 nsew
flabel metal1 819 1185 1019 1385 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal1 1809 1258 2009 1458 0 FreeSans 256 0 0 0 DGND
port 4 nsew
flabel metal1 1570 1249 1770 1449 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 825 -6 1025 194 0 FreeSans 256 0 0 0 IN3
port 5 nsew
flabel metal1 815 895 1015 1095 0 FreeSans 256 0 0 0 IN1
port 0 nsew
<< end >>
