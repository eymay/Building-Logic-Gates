** sch_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/xschem/NAND3/NAND3_eymenunay_TB.sch
**.subckt NAND3_eymenunay_TB
VDD VDD GND 1.8
V2 IN1 GND pulse 0 1.8 0n 1n 1n 100n 200n
V1 IN2 GND pulse 0 1.8 50n 1n 1n 100n 200n
X1 IN1 IN3 VDD GND OUT IN2 NAND3_eymenunay
V3 IN3 GND pulse 0 1.8 75n 1n 1n 100n 200n
C1 OUT GND 100f m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm




.control

tran 0.1n 400n
save all
plot IN1 IN2 IN3 OUT



.endc


**** end user architecture code
**.ends

* expanding   symbol:  NAND3_eymenunay.sym # of pins=6
** sym_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/xschem/NAND3/NAND3_eymenunay.sym
** sch_path: /home/ubuntu/Desktop/examples/xschem/VLSI-II/xschem/NAND3/NAND3_eymenunay.sch
.subckt NAND3_eymenunay  IN1 IN3 DVDD DGND OUT IN2
*.ipin IN1
*.ipin IN2
*.opin OUT
*.iopin DVDD
*.iopin DGND
*.ipin IN3
XM1 OUT IN1 net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 IN2 net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT IN1 DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT IN2 DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT IN3 DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 IN3 DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
